*** SPICE deck for cell mux{lay} from library gates_ma
*** Created on Thu Sep 26, 2013 07:43:08
*** Last revised on Fri Sep 27, 2013 14:42:50
*** Written on Fri Sep 27, 2013 14:47:25 by Electric VLSI Design System, 
*version 9.04
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

*** TOP LEVEL CELL: mux{lay}
Mnmos@5 gnd S net@228 gnd N L=0.6U W=1.2U AS=7.11P AD=5.4P PS=11.175U 
+PD=13.8U
Mnmos@6 net@222 D0 gnd gnd N L=0.6U W=1.2U AS=5.4P AD=1.8P PS=13.8U PD=4.2U
Mnmos@7 Yb net@228 net@222 gnd N L=0.6U W=1.2U AS=1.8P AD=5.22P PS=4.2U 
+PD=7.425U
Mnmos@8 net@225 S Yb gnd N L=0.6U W=1.2U AS=5.22P AD=1.62P PS=7.425U PD=3.9U
Mnmos@9 gnd D1 net@225 gnd N L=0.6U W=1.2U AS=1.62P AD=5.4P PS=3.9U PD=13.8U
Mpmos@0 vdd S net@228 vdd P L=0.6U W=2.4U AS=7.11P AD=10.26P PS=11.175U 
+PD=16.55U
Mpmos@1 net@215 D0 vdd vdd P L=0.6U W=2.4U AS=10.26P AD=4.14P PS=16.55U 
+PD=5.85U
Mpmos@2 Yb S net@215 vdd P L=0.6U W=2.4U AS=4.14P AD=5.22P PS=5.85U PD=7.425U
Mpmos@3 net@218 net@228 Yb vdd P L=0.6U W=2.4U AS=5.22P AD=4.14P PS=7.425U 
+PD=5.85U
Mpmos@4 vdd D1 net@218 vdd P L=0.6U W=2.4U AS=4.14P AD=10.26P PS=5.85U 
+PD=16.55U
.END
